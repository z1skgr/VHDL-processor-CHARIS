----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    00:31:07 02/22/2018 
-- Design Name: 
-- Module Name:    ALUSTAGE - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity ALUSTAGE is
    Port ( RF_A : in  STD_LOGIC_VECTOR (31 downto 0);
           RF_B : in  STD_LOGIC_VECTOR (31 downto 0);
           Immed : in  STD_LOGIC_VECTOR (31 downto 0);
           ALU_Bin_sel : in  STD_LOGIC;
			  ALU_Ain_sel : in  STD_LOGIC;
			  ALU_Cin_sel:in std_logic;
			  ALU_Din_sel:in std_logic;
			  ALU_Ein_sel:in std_logic;
			  ALU_func : in  STD_LOGIC_VECTOR (3 downto 0);
			  Zero:out std_logic;
           ALU_out : out  STD_LOGIC_VECTOR (31 downto 0));
end ALUSTAGE;

architecture Behavioral of ALUSTAGE is
component ALU is
    Port ( A : in  STD_LOGIC_VECTOR (31 downto 0);
           B : in  STD_LOGIC_VECTOR (31 downto 0);
           Op : in  STD_LOGIC_VECTOR (3 downto 0);
           Outp : out  STD_LOGIC_VECTOR (31 downto 0);
           Zero : out  STD_LOGIC;
           Cout : out  STD_LOGIC;
           Ovf : out  STD_LOGIC);
end component;

component Mux2to1_32bit is
	port(	Q0 : in  STD_LOGIC_VECTOR(31 downto 0);
         Q1 : in  STD_LOGIC_VECTOR(31 downto 0);
         Sign : in  STD_LOGIC;
         Outm : out  STD_LOGIC_VECTOR(31 downto 0));
end component;

signal mout5,mout4,mout3,mout1,mout2:STD_LOGIC_VECTOR(31 downto 0);

begin
ALUM:ALU
    port map(A=>mout1,
             B=>mout5,
             Op=>ALU_func,
				 Zero=>Zero,
             Outp =>ALU_out
	          );
Mux2:Mux2to1_32bit
      port map(Q0 =>RF_B,
               Q1 =>Immed,
               Sign =>ALU_Bin_sel,
               Outm =>mout2
		         );

Mux5:Mux2to1_32bit
      port map(Q0 =>mout2,
               Q1 =>"00000000000000000000000000000001",
               Sign =>ALU_Ein_sel,
               Outm =>mout5
		         );					

					
Mux1:Mux2to1_32bit
port map(Q0 =>RF_A,
               Q1 =>mout4,
               Sign =>ALU_Ain_sel,
               Outm =>mout1
		         );
					

Mux3:Mux2to1_32bit
port map(Q0=>"00000000000000000000000000000000",
			Q1=>RF_B,
			Sign=>ALU_Cin_sel,
			Outm=>mout3);
			
Mux4:Mux2to1_32bit
port map(Q0=>mout3,
			Q1=>"00000000000000000000000000000001",
			Sign=>ALU_Din_sel,
			Outm=>mout4
);

end Behavioral;

